`ifndef _global_vh_
`define _global_vh_

/**** Memory setup ****/
`define MEM_SIZE     'h10_0000

`define CHANNEL_SIZE    8
`define PIXEL_SIZE      24

/**** Input/output files ****/
`define IFILE       "imgs/red.bmp"
`define OFILE       "out/red_out.bmp"

/**** Testbench setup ****/
`define SIM_TIME 8_000_000

`endif
