`ifndef _global_vh_
`define _global_vh_

/**** Memory setup ****/
`define MEM_SIZE     'h10_0000

`define CHANNEL_SIZE    8
`define PIXEL_SIZE      24

/**** Input/output files ****/
`define IFILE       "imgs/balloon.bmp"
`define OFILE       "out/out.bmp"

/**** Testbench setup ****/
`define SIM_TIME 6_000_000

`endif
